//
// orpsoc-defines
//
`define MOR1KX
`define UART0
`define SPI0
`define JTAG_DEBUG
`define RAM_WB
`define BOOTROM
// end of included module defines - keep this comment line here
